// Clock generator module file
// frequencies -> 32f -> 4f -> 2f -> f
